
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom1 is
generic
	(
		ADDR_WIDTH : integer := 15 -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture rtl of controller_rom1 is

	signal addr1 : integer range 0 to 2**ADDR_WIDTH-1;

	--  build up 2D array to hold the memory
	type word_t is array (0 to 3) of std_logic_vector(7 downto 0);
	type ram_t is array (0 to 2 ** ADDR_WIDTH - 1) of word_t;

	signal ram : ram_t:=
	(

     0 => (x"04",x"87",x"da",x"01"),
     1 => (x"58",x"0e",x"87",x"dd"),
     2 => (x"0e",x"5a",x"59",x"5e"),
     3 => (x"00",x"00",x"29",x"27"),
     4 => (x"4a",x"26",x"0f",x"00"),
     5 => (x"48",x"26",x"49",x"26"),
     6 => (x"08",x"26",x"80",x"ff"),
     7 => (x"00",x"2d",x"27",x"4f"),
     8 => (x"27",x"4f",x"00",x"00"),
     9 => (x"00",x"00",x"00",x"2a"),
    10 => (x"fd",x"00",x"4f",x"4f"),
    11 => (x"dc",x"d0",x"c1",x"87"),
    12 => (x"48",x"c0",x"c8",x"4e"),
    13 => (x"d5",x"c1",x"28",x"c2"),
    14 => (x"ea",x"d6",x"e5",x"ea"),
    15 => (x"c1",x"46",x"71",x"49"),
    16 => (x"87",x"f9",x"01",x"88"),
    17 => (x"49",x"dc",x"d0",x"c1"),
    18 => (x"48",x"d0",x"cc",x"c1"),
    19 => (x"03",x"89",x"d0",x"89"),
    20 => (x"40",x"40",x"40",x"c0"),
    21 => (x"d0",x"87",x"f6",x"40"),
    22 => (x"50",x"c0",x"05",x"81"),
    23 => (x"f9",x"05",x"89",x"c1"),
    24 => (x"cd",x"cc",x"c1",x"87"),
    25 => (x"c9",x"cc",x"c1",x"4d"),
    26 => (x"02",x"ad",x"74",x"4c"),
    27 => (x"0f",x"24",x"87",x"c4"),
    28 => (x"c2",x"dc",x"87",x"f7"),
    29 => (x"cd",x"cc",x"c1",x"87"),
    30 => (x"cd",x"cc",x"c1",x"4d"),
    31 => (x"02",x"ad",x"74",x"4c"),
    32 => (x"8c",x"c4",x"87",x"c6"),
    33 => (x"87",x"f5",x"0f",x"6c"),
    34 => (x"1e",x"87",x"fd",x"00"),
    35 => (x"4a",x"71",x"86",x"fc"),
    36 => (x"69",x"49",x"c0",x"ff"),
    37 => (x"98",x"c0",x"c4",x"48"),
    38 => (x"98",x"48",x"7e",x"70"),
    39 => (x"72",x"87",x"f4",x"02"),
    40 => (x"8e",x"fc",x"48",x"79"),
    41 => (x"73",x"1e",x"4f",x"26"),
    42 => (x"a9",x"73",x"81",x"48"),
    43 => (x"12",x"87",x"c5",x"02"),
    44 => (x"87",x"f6",x"05",x"53"),
    45 => (x"ff",x"1e",x"4f",x"26"),
    46 => (x"ff",x"c3",x"48",x"d4"),
    47 => (x"26",x"48",x"68",x"78"),
    48 => (x"d4",x"ff",x"1e",x"4f"),
    49 => (x"78",x"ff",x"c3",x"48"),
    50 => (x"c0",x"48",x"d0",x"ff"),
    51 => (x"d4",x"ff",x"78",x"e1"),
    52 => (x"26",x"78",x"d4",x"48"),
    53 => (x"d0",x"ff",x"1e",x"4f"),
    54 => (x"78",x"e0",x"c0",x"48"),
    55 => (x"ff",x"1e",x"4f",x"26"),
    56 => (x"49",x"70",x"87",x"d4"),
    57 => (x"87",x"c6",x"02",x"99"),
    58 => (x"05",x"a9",x"fb",x"c0"),
    59 => (x"48",x"71",x"87",x"f1"),
    60 => (x"5e",x"0e",x"4f",x"26"),
    61 => (x"71",x"0e",x"5c",x"5b"),
    62 => (x"fe",x"4c",x"c0",x"4b"),
    63 => (x"49",x"70",x"87",x"f8"),
    64 => (x"f9",x"c0",x"02",x"99"),
    65 => (x"a9",x"ec",x"c0",x"87"),
    66 => (x"87",x"f2",x"c0",x"02"),
    67 => (x"02",x"a9",x"fb",x"c0"),
    68 => (x"cc",x"87",x"eb",x"c0"),
    69 => (x"03",x"ac",x"b7",x"66"),
    70 => (x"66",x"d0",x"87",x"c7"),
    71 => (x"71",x"87",x"c2",x"02"),
    72 => (x"02",x"99",x"71",x"53"),
    73 => (x"84",x"c1",x"87",x"c2"),
    74 => (x"70",x"87",x"cb",x"fe"),
    75 => (x"cd",x"02",x"99",x"49"),
    76 => (x"a9",x"ec",x"c0",x"87"),
    77 => (x"c0",x"87",x"c7",x"02"),
    78 => (x"ff",x"05",x"a9",x"fb"),
    79 => (x"66",x"d0",x"87",x"d5"),
    80 => (x"c0",x"87",x"c3",x"02"),
    81 => (x"ec",x"c0",x"7b",x"97"),
    82 => (x"87",x"c4",x"05",x"a9"),
    83 => (x"87",x"c5",x"4a",x"74"),
    84 => (x"0a",x"c0",x"4a",x"74"),
    85 => (x"26",x"48",x"72",x"8a"),
    86 => (x"26",x"4b",x"26",x"4c"),
    87 => (x"d5",x"fd",x"1e",x"4f"),
    88 => (x"4a",x"49",x"70",x"87"),
    89 => (x"04",x"aa",x"f0",x"c0"),
    90 => (x"f9",x"c0",x"87",x"c9"),
    91 => (x"87",x"c3",x"01",x"aa"),
    92 => (x"c1",x"8a",x"f0",x"c0"),
    93 => (x"c9",x"04",x"aa",x"c1"),
    94 => (x"aa",x"da",x"c1",x"87"),
    95 => (x"c0",x"87",x"c3",x"01"),
    96 => (x"48",x"72",x"8a",x"f7"),
    97 => (x"26",x"1e",x"4f",x"26"),
    98 => (x"4f",x"26",x"1e",x"4f"),
    99 => (x"1e",x"4f",x"26",x"1e"),
   100 => (x"f7",x"c0",x"49",x"c0"),
   101 => (x"4f",x"26",x"87",x"ef"),
   102 => (x"49",x"4a",x"71",x"1e"),
   103 => (x"dc",x"df",x"91",x"cc"),
   104 => (x"c1",x"81",x"c8",x"81"),
   105 => (x"11",x"48",x"d4",x"cc"),
   106 => (x"a2",x"f0",x"c0",x"50"),
   107 => (x"87",x"db",x"fb",x"49"),
   108 => (x"de",x"d6",x"49",x"c0"),
   109 => (x"1e",x"4f",x"26",x"87"),
   110 => (x"c3",x"4a",x"d4",x"ff"),
   111 => (x"d0",x"ff",x"7a",x"ff"),
   112 => (x"78",x"e1",x"c0",x"48"),
   113 => (x"7a",x"71",x"7a",x"de"),
   114 => (x"28",x"b7",x"c8",x"48"),
   115 => (x"48",x"71",x"7a",x"70"),
   116 => (x"70",x"28",x"b7",x"d0"),
   117 => (x"d8",x"48",x"71",x"7a"),
   118 => (x"7a",x"70",x"28",x"b7"),
   119 => (x"c0",x"48",x"d0",x"ff"),
   120 => (x"4f",x"26",x"78",x"e0"),
   121 => (x"5c",x"5b",x"5e",x"0e"),
   122 => (x"86",x"f4",x"0e",x"5d"),
   123 => (x"cc",x"49",x"4d",x"71"),
   124 => (x"81",x"dc",x"df",x"91"),
   125 => (x"ca",x"4a",x"a1",x"c8"),
   126 => (x"a6",x"c4",x"7e",x"a1"),
   127 => (x"d0",x"cc",x"c1",x"48"),
   128 => (x"97",x"6e",x"78",x"bf"),
   129 => (x"66",x"c4",x"4b",x"bf"),
   130 => (x"12",x"2c",x"73",x"4c"),
   131 => (x"58",x"a6",x"cc",x"48"),
   132 => (x"84",x"c1",x"9c",x"70"),
   133 => (x"69",x"97",x"81",x"c9"),
   134 => (x"04",x"ac",x"b7",x"49"),
   135 => (x"4c",x"c0",x"87",x"c2"),
   136 => (x"4a",x"bf",x"97",x"6e"),
   137 => (x"72",x"49",x"66",x"c8"),
   138 => (x"c4",x"b9",x"ff",x"31"),
   139 => (x"48",x"74",x"99",x"66"),
   140 => (x"4a",x"70",x"30",x"72"),
   141 => (x"d4",x"cc",x"c1",x"b1"),
   142 => (x"fa",x"fd",x"71",x"59"),
   143 => (x"c1",x"1e",x"c7",x"87"),
   144 => (x"1e",x"bf",x"d8",x"cc"),
   145 => (x"c1",x"1e",x"dc",x"df"),
   146 => (x"bf",x"97",x"d4",x"cc"),
   147 => (x"87",x"f3",x"c1",x"49"),
   148 => (x"f3",x"c0",x"49",x"75"),
   149 => (x"8e",x"e8",x"87",x"ce"),
   150 => (x"4c",x"26",x"4d",x"26"),
   151 => (x"4f",x"26",x"4b",x"26"),
   152 => (x"71",x"1e",x"73",x"1e"),
   153 => (x"fb",x"fd",x"49",x"4b"),
   154 => (x"fd",x"49",x"73",x"87"),
   155 => (x"4b",x"26",x"87",x"f6"),
   156 => (x"73",x"1e",x"4f",x"26"),
   157 => (x"c2",x"4b",x"71",x"1e"),
   158 => (x"d6",x"02",x"4a",x"a3"),
   159 => (x"05",x"8a",x"c1",x"87"),
   160 => (x"c1",x"87",x"e2",x"c0"),
   161 => (x"02",x"bf",x"d8",x"cc"),
   162 => (x"c1",x"48",x"87",x"db"),
   163 => (x"dc",x"cc",x"c1",x"88"),
   164 => (x"c1",x"87",x"d2",x"58"),
   165 => (x"02",x"bf",x"dc",x"cc"),
   166 => (x"cc",x"c1",x"87",x"cb"),
   167 => (x"c1",x"48",x"bf",x"d8"),
   168 => (x"dc",x"cc",x"c1",x"80"),
   169 => (x"c1",x"1e",x"c7",x"58"),
   170 => (x"1e",x"bf",x"d8",x"cc"),
   171 => (x"c1",x"1e",x"dc",x"df"),
   172 => (x"bf",x"97",x"d4",x"cc"),
   173 => (x"73",x"87",x"cc",x"49"),
   174 => (x"e7",x"f1",x"c0",x"49"),
   175 => (x"26",x"8e",x"f4",x"87"),
   176 => (x"0e",x"4f",x"26",x"4b"),
   177 => (x"5d",x"5c",x"5b",x"5e"),
   178 => (x"86",x"cc",x"ff",x"0e"),
   179 => (x"59",x"a6",x"e4",x"c0"),
   180 => (x"c0",x"48",x"a6",x"cc"),
   181 => (x"c0",x"80",x"c4",x"78"),
   182 => (x"c1",x"80",x"c4",x"78"),
   183 => (x"c4",x"78",x"66",x"c8"),
   184 => (x"c4",x"78",x"c1",x"80"),
   185 => (x"c1",x"78",x"c1",x"80"),
   186 => (x"c1",x"48",x"dc",x"cc"),
   187 => (x"87",x"d1",x"f7",x"78"),
   188 => (x"f7",x"87",x"eb",x"f7"),
   189 => (x"4c",x"70",x"87",x"c0"),
   190 => (x"02",x"ac",x"fb",x"c0"),
   191 => (x"c0",x"87",x"ef",x"c1"),
   192 => (x"c1",x"05",x"66",x"e0"),
   193 => (x"c4",x"c1",x"87",x"e5"),
   194 => (x"82",x"c4",x"4a",x"66"),
   195 => (x"f4",x"dc",x"7e",x"6a"),
   196 => (x"20",x"49",x"6e",x"48"),
   197 => (x"10",x"41",x"20",x"41"),
   198 => (x"66",x"c4",x"c1",x"51"),
   199 => (x"78",x"c6",x"c6",x"48"),
   200 => (x"81",x"c7",x"49",x"6a"),
   201 => (x"c4",x"c1",x"51",x"74"),
   202 => (x"81",x"c8",x"49",x"66"),
   203 => (x"a6",x"d8",x"51",x"c1"),
   204 => (x"c1",x"78",x"c2",x"48"),
   205 => (x"c9",x"49",x"66",x"c4"),
   206 => (x"c1",x"51",x"c0",x"81"),
   207 => (x"ca",x"49",x"66",x"c4"),
   208 => (x"c1",x"51",x"c0",x"81"),
   209 => (x"6a",x"1e",x"d8",x"1e"),
   210 => (x"f6",x"81",x"c8",x"49"),
   211 => (x"86",x"c8",x"87",x"e4"),
   212 => (x"48",x"66",x"c8",x"c1"),
   213 => (x"c7",x"01",x"a8",x"c0"),
   214 => (x"48",x"a6",x"d0",x"87"),
   215 => (x"87",x"ce",x"78",x"c1"),
   216 => (x"48",x"66",x"c8",x"c1"),
   217 => (x"a6",x"d8",x"88",x"c1"),
   218 => (x"f5",x"87",x"c3",x"58"),
   219 => (x"9c",x"74",x"87",x"f0"),
   220 => (x"87",x"c0",x"cd",x"02"),
   221 => (x"c1",x"48",x"66",x"d0"),
   222 => (x"03",x"a8",x"66",x"cc"),
   223 => (x"c8",x"87",x"f5",x"cc"),
   224 => (x"78",x"c0",x"48",x"a6"),
   225 => (x"87",x"ee",x"f4",x"7e"),
   226 => (x"d0",x"c1",x"4c",x"70"),
   227 => (x"e2",x"c2",x"05",x"ac"),
   228 => (x"48",x"a6",x"c4",x"87"),
   229 => (x"c4",x"f7",x"78",x"6e"),
   230 => (x"48",x"7e",x"70",x"87"),
   231 => (x"06",x"a8",x"66",x"cc"),
   232 => (x"a6",x"cc",x"87",x"c5"),
   233 => (x"f4",x"78",x"6e",x"48"),
   234 => (x"4c",x"70",x"87",x"cc"),
   235 => (x"05",x"ac",x"ec",x"c0"),
   236 => (x"d0",x"87",x"ea",x"c1"),
   237 => (x"91",x"cc",x"49",x"66"),
   238 => (x"81",x"66",x"c4",x"c1"),
   239 => (x"6a",x"4a",x"a1",x"c4"),
   240 => (x"4a",x"a1",x"c8",x"4d"),
   241 => (x"d8",x"c6",x"52",x"6e"),
   242 => (x"87",x"ea",x"f3",x"79"),
   243 => (x"02",x"9c",x"4c",x"70"),
   244 => (x"fb",x"c0",x"87",x"d8"),
   245 => (x"87",x"d2",x"02",x"ac"),
   246 => (x"d9",x"f3",x"55",x"74"),
   247 => (x"9c",x"4c",x"70",x"87"),
   248 => (x"c0",x"87",x"c7",x"02"),
   249 => (x"ff",x"05",x"ac",x"fb"),
   250 => (x"e0",x"c0",x"87",x"ee"),
   251 => (x"55",x"c1",x"c2",x"55"),
   252 => (x"c0",x"7d",x"97",x"c0"),
   253 => (x"c4",x"48",x"66",x"e0"),
   254 => (x"db",x"05",x"a8",x"66"),
   255 => (x"48",x"66",x"d0",x"87"),
   256 => (x"04",x"a8",x"66",x"d4"),
   257 => (x"66",x"d0",x"87",x"ca"),
   258 => (x"d4",x"80",x"c1",x"48"),
   259 => (x"87",x"c8",x"58",x"a6"),
   260 => (x"c1",x"48",x"66",x"d4"),
   261 => (x"58",x"a6",x"d8",x"88"),
   262 => (x"70",x"87",x"db",x"f2"),
   263 => (x"ac",x"d0",x"c1",x"4c"),
   264 => (x"dc",x"87",x"c9",x"05"),
   265 => (x"80",x"c1",x"48",x"66"),
   266 => (x"58",x"a6",x"e0",x"c0"),
   267 => (x"02",x"ac",x"d0",x"c1"),
   268 => (x"6e",x"87",x"de",x"fd"),
   269 => (x"66",x"e0",x"c0",x"48"),
   270 => (x"d8",x"c9",x"05",x"a8"),
   271 => (x"a6",x"e4",x"c0",x"87"),
   272 => (x"74",x"78",x"c0",x"48"),
   273 => (x"88",x"fb",x"c0",x"48"),
   274 => (x"70",x"58",x"a6",x"c8"),
   275 => (x"c9",x"c9",x"02",x"98"),
   276 => (x"88",x"cb",x"48",x"87"),
   277 => (x"70",x"58",x"a6",x"c8"),
   278 => (x"cc",x"c1",x"02",x"98"),
   279 => (x"88",x"c9",x"48",x"87"),
   280 => (x"70",x"58",x"a6",x"c8"),
   281 => (x"f6",x"c3",x"02",x"98"),
   282 => (x"88",x"c4",x"48",x"87"),
   283 => (x"70",x"58",x"a6",x"c8"),
   284 => (x"87",x"cf",x"02",x"98"),
   285 => (x"c8",x"88",x"c1",x"48"),
   286 => (x"98",x"70",x"58",x"a6"),
   287 => (x"87",x"df",x"c3",x"02"),
   288 => (x"c8",x"87",x"ca",x"c8"),
   289 => (x"f0",x"c0",x"48",x"a6"),
   290 => (x"87",x"ea",x"f0",x"78"),
   291 => (x"ec",x"c0",x"4c",x"70"),
   292 => (x"87",x"c3",x"02",x"ac"),
   293 => (x"c0",x"5c",x"a6",x"cc"),
   294 => (x"cc",x"02",x"ac",x"ec"),
   295 => (x"87",x"d6",x"f0",x"87"),
   296 => (x"ec",x"c0",x"4c",x"70"),
   297 => (x"f4",x"ff",x"05",x"ac"),
   298 => (x"ac",x"ec",x"c0",x"87"),
   299 => (x"f0",x"87",x"c3",x"02"),
   300 => (x"1e",x"c0",x"87",x"c4"),
   301 => (x"66",x"d8",x"1e",x"ca"),
   302 => (x"c1",x"91",x"cc",x"49"),
   303 => (x"71",x"48",x"66",x"cc"),
   304 => (x"58",x"a6",x"cc",x"80"),
   305 => (x"c4",x"48",x"66",x"c8"),
   306 => (x"58",x"a6",x"d0",x"80"),
   307 => (x"49",x"bf",x"66",x"cc"),
   308 => (x"c1",x"87",x"df",x"f0"),
   309 => (x"d4",x"1e",x"de",x"1e"),
   310 => (x"f0",x"49",x"bf",x"66"),
   311 => (x"86",x"d0",x"87",x"d4"),
   312 => (x"c0",x"48",x"49",x"70"),
   313 => (x"ec",x"c0",x"88",x"08"),
   314 => (x"a8",x"c0",x"58",x"a6"),
   315 => (x"87",x"ee",x"c0",x"06"),
   316 => (x"48",x"66",x"e8",x"c0"),
   317 => (x"c0",x"03",x"a8",x"dd"),
   318 => (x"66",x"c4",x"87",x"e4"),
   319 => (x"e8",x"c0",x"49",x"bf"),
   320 => (x"e0",x"c0",x"81",x"66"),
   321 => (x"66",x"e8",x"c0",x"51"),
   322 => (x"c4",x"81",x"c1",x"49"),
   323 => (x"c2",x"81",x"bf",x"66"),
   324 => (x"e8",x"c0",x"51",x"c1"),
   325 => (x"81",x"c2",x"49",x"66"),
   326 => (x"81",x"bf",x"66",x"c4"),
   327 => (x"48",x"6e",x"51",x"c0"),
   328 => (x"6e",x"78",x"c6",x"c6"),
   329 => (x"d8",x"81",x"c8",x"49"),
   330 => (x"49",x"6e",x"51",x"66"),
   331 => (x"66",x"dc",x"81",x"c9"),
   332 => (x"ca",x"49",x"6e",x"51"),
   333 => (x"51",x"66",x"c8",x"81"),
   334 => (x"c1",x"48",x"66",x"d8"),
   335 => (x"58",x"a6",x"dc",x"80"),
   336 => (x"d4",x"48",x"66",x"d0"),
   337 => (x"cb",x"04",x"a8",x"66"),
   338 => (x"48",x"66",x"d0",x"87"),
   339 => (x"a6",x"d4",x"80",x"c1"),
   340 => (x"87",x"c6",x"c5",x"58"),
   341 => (x"c1",x"48",x"66",x"d4"),
   342 => (x"58",x"a6",x"d8",x"88"),
   343 => (x"ef",x"87",x"fb",x"c4"),
   344 => (x"ec",x"c0",x"87",x"fb"),
   345 => (x"f4",x"ef",x"58",x"a6"),
   346 => (x"a6",x"f0",x"c0",x"87"),
   347 => (x"a8",x"ec",x"c0",x"58"),
   348 => (x"87",x"c9",x"c0",x"05"),
   349 => (x"e8",x"c0",x"48",x"a6"),
   350 => (x"c3",x"c0",x"78",x"66"),
   351 => (x"87",x"f6",x"ec",x"87"),
   352 => (x"cc",x"49",x"66",x"d0"),
   353 => (x"66",x"c4",x"c1",x"91"),
   354 => (x"c8",x"80",x"71",x"48"),
   355 => (x"66",x"c4",x"58",x"a6"),
   356 => (x"c4",x"82",x"c8",x"4a"),
   357 => (x"81",x"ca",x"49",x"66"),
   358 => (x"51",x"66",x"e8",x"c0"),
   359 => (x"49",x"66",x"ec",x"c0"),
   360 => (x"e8",x"c0",x"81",x"c1"),
   361 => (x"48",x"c1",x"89",x"66"),
   362 => (x"49",x"70",x"30",x"71"),
   363 => (x"97",x"71",x"89",x"c1"),
   364 => (x"d0",x"cc",x"c1",x"7a"),
   365 => (x"e8",x"c0",x"49",x"bf"),
   366 => (x"6a",x"97",x"29",x"66"),
   367 => (x"98",x"71",x"48",x"4a"),
   368 => (x"58",x"a6",x"f4",x"c0"),
   369 => (x"c4",x"48",x"66",x"c4"),
   370 => (x"58",x"a6",x"cc",x"80"),
   371 => (x"4d",x"bf",x"66",x"c8"),
   372 => (x"48",x"66",x"e0",x"c0"),
   373 => (x"c0",x"02",x"a8",x"6e"),
   374 => (x"7e",x"c0",x"87",x"c5"),
   375 => (x"c1",x"87",x"c2",x"c0"),
   376 => (x"c0",x"1e",x"6e",x"7e"),
   377 => (x"49",x"75",x"1e",x"e0"),
   378 => (x"c8",x"87",x"c7",x"ec"),
   379 => (x"c0",x"4c",x"70",x"86"),
   380 => (x"c1",x"06",x"ac",x"b7"),
   381 => (x"85",x"74",x"87",x"d1"),
   382 => (x"49",x"bf",x"66",x"c8"),
   383 => (x"75",x"81",x"e0",x"c0"),
   384 => (x"c0",x"dd",x"4b",x"89"),
   385 => (x"dd",x"ea",x"71",x"4a"),
   386 => (x"75",x"85",x"c2",x"87"),
   387 => (x"66",x"e4",x"c0",x"7e"),
   388 => (x"c0",x"80",x"c1",x"48"),
   389 => (x"c0",x"58",x"a6",x"e8"),
   390 => (x"c1",x"49",x"66",x"f0"),
   391 => (x"02",x"a9",x"70",x"81"),
   392 => (x"c0",x"87",x"c5",x"c0"),
   393 => (x"87",x"c2",x"c0",x"4d"),
   394 => (x"1e",x"75",x"4d",x"c1"),
   395 => (x"49",x"bf",x"66",x"cc"),
   396 => (x"c4",x"81",x"e0",x"c0"),
   397 => (x"1e",x"71",x"89",x"66"),
   398 => (x"ea",x"49",x"66",x"c8"),
   399 => (x"86",x"c8",x"87",x"f4"),
   400 => (x"01",x"a8",x"b7",x"c0"),
   401 => (x"c0",x"87",x"c6",x"ff"),
   402 => (x"c0",x"02",x"66",x"e4"),
   403 => (x"66",x"c4",x"87",x"d2"),
   404 => (x"c0",x"81",x"c9",x"49"),
   405 => (x"c4",x"51",x"66",x"e4"),
   406 => (x"e4",x"c7",x"48",x"66"),
   407 => (x"87",x"cd",x"c0",x"78"),
   408 => (x"c9",x"49",x"66",x"c4"),
   409 => (x"c4",x"51",x"c2",x"81"),
   410 => (x"e0",x"c9",x"48",x"66"),
   411 => (x"48",x"66",x"d0",x"78"),
   412 => (x"04",x"a8",x"66",x"d4"),
   413 => (x"d0",x"87",x"cb",x"c0"),
   414 => (x"80",x"c1",x"48",x"66"),
   415 => (x"c0",x"58",x"a6",x"d4"),
   416 => (x"66",x"d4",x"87",x"d8"),
   417 => (x"d8",x"88",x"c1",x"48"),
   418 => (x"cd",x"c0",x"58",x"a6"),
   419 => (x"87",x"ce",x"e9",x"87"),
   420 => (x"c5",x"c0",x"4c",x"70"),
   421 => (x"87",x"c6",x"e9",x"87"),
   422 => (x"66",x"dc",x"4c",x"70"),
   423 => (x"c0",x"80",x"c1",x"48"),
   424 => (x"74",x"58",x"a6",x"e0"),
   425 => (x"cb",x"c0",x"02",x"9c"),
   426 => (x"48",x"66",x"d0",x"87"),
   427 => (x"a8",x"66",x"cc",x"c1"),
   428 => (x"87",x"cb",x"f3",x"04"),
   429 => (x"c7",x"48",x"66",x"d0"),
   430 => (x"e1",x"c0",x"03",x"a8"),
   431 => (x"4c",x"66",x"d0",x"87"),
   432 => (x"48",x"dc",x"cc",x"c1"),
   433 => (x"49",x"74",x"78",x"c0"),
   434 => (x"c4",x"c1",x"91",x"cc"),
   435 => (x"a1",x"c4",x"81",x"66"),
   436 => (x"c0",x"4a",x"6a",x"4a"),
   437 => (x"84",x"c1",x"79",x"52"),
   438 => (x"ff",x"04",x"ac",x"c7"),
   439 => (x"e0",x"c0",x"87",x"e2"),
   440 => (x"e0",x"c0",x"02",x"66"),
   441 => (x"66",x"c4",x"c1",x"87"),
   442 => (x"81",x"d4",x"c1",x"49"),
   443 => (x"4a",x"66",x"c4",x"c1"),
   444 => (x"c0",x"82",x"dc",x"c1"),
   445 => (x"79",x"d8",x"c6",x"52"),
   446 => (x"49",x"66",x"c4",x"c1"),
   447 => (x"dd",x"81",x"d8",x"c1"),
   448 => (x"d4",x"c0",x"79",x"c4"),
   449 => (x"66",x"c4",x"c1",x"87"),
   450 => (x"81",x"d4",x"c1",x"49"),
   451 => (x"4a",x"66",x"c4",x"c1"),
   452 => (x"dd",x"82",x"d8",x"c1"),
   453 => (x"cf",x"c6",x"7a",x"cc"),
   454 => (x"66",x"c4",x"c1",x"79"),
   455 => (x"81",x"e0",x"c1",x"49"),
   456 => (x"e6",x"79",x"f2",x"c9"),
   457 => (x"66",x"cc",x"87",x"ef"),
   458 => (x"8e",x"cc",x"ff",x"48"),
   459 => (x"4c",x"26",x"4d",x"26"),
   460 => (x"4f",x"26",x"4b",x"26"),
   461 => (x"64",x"61",x"6f",x"4c"),
   462 => (x"20",x"2e",x"2a",x"20"),
   463 => (x"00",x"00",x"00",x"00"),
   464 => (x"00",x"00",x"20",x"3a"),
   465 => (x"61",x"42",x"20",x"80"),
   466 => (x"00",x"00",x"6b",x"63"),
   467 => (x"78",x"45",x"20",x"80"),
   468 => (x"1e",x"00",x"74",x"69"),
   469 => (x"cc",x"c1",x"1e",x"c7"),
   470 => (x"df",x"1e",x"bf",x"d8"),
   471 => (x"cc",x"c1",x"1e",x"dc"),
   472 => (x"49",x"bf",x"97",x"d4"),
   473 => (x"df",x"87",x"dc",x"ed"),
   474 => (x"e0",x"c0",x"49",x"dc"),
   475 => (x"8e",x"f4",x"87",x"c4"),
   476 => (x"c0",x"1e",x"4f",x"26"),
   477 => (x"1e",x"4f",x"26",x"48"),
   478 => (x"c0",x"87",x"fa",x"c6"),
   479 => (x"df",x"48",x"f4",x"e0"),
   480 => (x"e8",x"fe",x"78",x"d0"),
   481 => (x"e9",x"df",x"49",x"a0"),
   482 => (x"de",x"49",x"c7",x"87"),
   483 => (x"49",x"c1",x"87",x"d6"),
   484 => (x"ff",x"87",x"f2",x"df"),
   485 => (x"ff",x"c3",x"48",x"d4"),
   486 => (x"d8",x"cc",x"c1",x"78"),
   487 => (x"c1",x"78",x"c0",x"48"),
   488 => (x"c0",x"48",x"d4",x"cc"),
   489 => (x"ea",x"fe",x"49",x"50"),
   490 => (x"87",x"c6",x"ff",x"87"),
   491 => (x"02",x"9a",x"4a",x"70"),
   492 => (x"e0",x"c0",x"87",x"cb"),
   493 => (x"49",x"c7",x"5a",x"f8"),
   494 => (x"c5",x"87",x"e9",x"dd"),
   495 => (x"df",x"49",x"c0",x"87"),
   496 => (x"ea",x"c2",x"87",x"c3"),
   497 => (x"e4",x"e0",x"c0",x"87"),
   498 => (x"26",x"87",x"fa",x"87"),
   499 => (x"00",x"00",x"00",x"4f"),
   500 => (x"74",x"6f",x"6f",x"42"),
   501 => (x"2e",x"67",x"6e",x"69"),
   502 => (x"00",x"00",x"2e",x"2e"),
   503 => (x"00",x"00",x"01",x"89"),
   504 => (x"00",x"00",x"13",x"20"),
   505 => (x"00",x"00",x"00",x"00"),
   506 => (x"00",x"00",x"01",x"89"),
   507 => (x"00",x"00",x"13",x"3e"),
   508 => (x"00",x"00",x"00",x"00"),
   509 => (x"00",x"00",x"01",x"89"),
   510 => (x"00",x"00",x"13",x"5c"),
   511 => (x"00",x"00",x"00",x"00"),
   512 => (x"00",x"00",x"01",x"89"),
   513 => (x"00",x"00",x"13",x"7a"),
   514 => (x"00",x"00",x"00",x"00"),
   515 => (x"00",x"00",x"01",x"89"),
   516 => (x"00",x"00",x"13",x"98"),
   517 => (x"00",x"00",x"00",x"00"),
   518 => (x"00",x"00",x"01",x"89"),
   519 => (x"00",x"00",x"13",x"b6"),
   520 => (x"00",x"00",x"00",x"00"),
   521 => (x"00",x"00",x"01",x"89"),
   522 => (x"00",x"00",x"13",x"d4"),
   523 => (x"00",x"00",x"00",x"00"),
   524 => (x"00",x"00",x"01",x"98"),
   525 => (x"00",x"00",x"00",x"00"),
   526 => (x"00",x"00",x"00",x"00"),
   527 => (x"00",x"00",x"01",x"8c"),
   528 => (x"00",x"00",x"00",x"00"),
   529 => (x"00",x"00",x"00",x"00"),
   530 => (x"db",x"86",x"fc",x"1e"),
   531 => (x"fc",x"7e",x"70",x"87"),
   532 => (x"1e",x"4f",x"26",x"8e"),
   533 => (x"c0",x"48",x"f0",x"fe"),
   534 => (x"79",x"09",x"cd",x"78"),
   535 => (x"1e",x"4f",x"26",x"09"),
   536 => (x"49",x"c8",x"e1",x"c0"),
   537 => (x"4f",x"26",x"87",x"ed"),
   538 => (x"bf",x"f0",x"fe",x"1e"),
   539 => (x"1e",x"4f",x"26",x"48"),
   540 => (x"c1",x"48",x"f0",x"fe"),
   541 => (x"1e",x"4f",x"26",x"78"),
   542 => (x"c0",x"48",x"f0",x"fe"),
   543 => (x"1e",x"4f",x"26",x"78"),
   544 => (x"52",x"c0",x"4a",x"71"),
   545 => (x"0e",x"4f",x"26",x"51"),
   546 => (x"5d",x"5c",x"5b",x"5e"),
   547 => (x"71",x"86",x"f4",x"0e"),
   548 => (x"7e",x"6d",x"97",x"4d"),
   549 => (x"97",x"4c",x"a5",x"c1"),
   550 => (x"a6",x"c8",x"48",x"6c"),
   551 => (x"c4",x"48",x"6e",x"58"),
   552 => (x"c5",x"05",x"a8",x"66"),
   553 => (x"c0",x"48",x"ff",x"87"),
   554 => (x"ca",x"ff",x"87",x"e6"),
   555 => (x"49",x"a5",x"c2",x"87"),
   556 => (x"71",x"4b",x"6c",x"97"),
   557 => (x"6b",x"97",x"4b",x"a3"),
   558 => (x"7e",x"6c",x"97",x"4b"),
   559 => (x"80",x"c1",x"48",x"6e"),
   560 => (x"c7",x"58",x"a6",x"c8"),
   561 => (x"58",x"a6",x"cc",x"98"),
   562 => (x"fe",x"7c",x"97",x"70"),
   563 => (x"48",x"73",x"87",x"e1"),
   564 => (x"4d",x"26",x"8e",x"f4"),
   565 => (x"4b",x"26",x"4c",x"26"),
   566 => (x"5e",x"0e",x"4f",x"26"),
   567 => (x"f4",x"0e",x"5c",x"5b"),
   568 => (x"d8",x"4c",x"71",x"86"),
   569 => (x"ff",x"c3",x"4a",x"66"),
   570 => (x"4b",x"a4",x"c2",x"9a"),
   571 => (x"73",x"49",x"6c",x"97"),
   572 => (x"51",x"72",x"49",x"a1"),
   573 => (x"6e",x"7e",x"6c",x"97"),
   574 => (x"c8",x"80",x"c1",x"48"),
   575 => (x"98",x"c7",x"58",x"a6"),
   576 => (x"70",x"58",x"a6",x"cc"),
   577 => (x"26",x"8e",x"f4",x"54"),
   578 => (x"26",x"4b",x"26",x"4c"),
   579 => (x"86",x"fc",x"1e",x"4f"),
   580 => (x"e0",x"87",x"e4",x"fd"),
   581 => (x"c0",x"49",x"4a",x"bf"),
   582 => (x"02",x"99",x"c0",x"e0"),
   583 => (x"1e",x"72",x"87",x"cb"),
   584 => (x"49",x"f4",x"cf",x"c1"),
   585 => (x"c4",x"87",x"f3",x"fe"),
   586 => (x"87",x"fc",x"fc",x"86"),
   587 => (x"fe",x"fc",x"7e",x"70"),
   588 => (x"26",x"8e",x"fc",x"87"),
   589 => (x"cf",x"c1",x"1e",x"4f"),
   590 => (x"c2",x"fd",x"49",x"f4"),
   591 => (x"cd",x"e4",x"c0",x"87"),
   592 => (x"87",x"cf",x"fc",x"49"),
   593 => (x"26",x"87",x"f1",x"c2"),
   594 => (x"1e",x"73",x"1e",x"4f"),
   595 => (x"49",x"f4",x"cf",x"c1"),
   596 => (x"70",x"87",x"f4",x"fc"),
   597 => (x"aa",x"b7",x"c0",x"4a"),
   598 => (x"87",x"cc",x"c2",x"04"),
   599 => (x"05",x"aa",x"f0",x"c3"),
   600 => (x"e7",x"c0",x"87",x"c9"),
   601 => (x"78",x"c1",x"48",x"f0"),
   602 => (x"c3",x"87",x"ed",x"c1"),
   603 => (x"c9",x"05",x"aa",x"e0"),
   604 => (x"f4",x"e7",x"c0",x"87"),
   605 => (x"c1",x"78",x"c1",x"48"),
   606 => (x"e7",x"c0",x"87",x"de"),
   607 => (x"c6",x"02",x"bf",x"f4"),
   608 => (x"a2",x"c0",x"c2",x"87"),
   609 => (x"72",x"87",x"c2",x"4b"),
   610 => (x"f0",x"e7",x"c0",x"4b"),
   611 => (x"e0",x"c0",x"02",x"bf"),
   612 => (x"c4",x"49",x"73",x"87"),
   613 => (x"c0",x"91",x"29",x"b7"),
   614 => (x"73",x"81",x"cc",x"e9"),
   615 => (x"c2",x"9a",x"cf",x"4a"),
   616 => (x"72",x"48",x"c1",x"92"),
   617 => (x"ff",x"4a",x"70",x"30"),
   618 => (x"69",x"48",x"72",x"ba"),
   619 => (x"db",x"79",x"70",x"98"),
   620 => (x"c4",x"49",x"73",x"87"),
   621 => (x"c0",x"91",x"29",x"b7"),
   622 => (x"73",x"81",x"cc",x"e9"),
   623 => (x"c2",x"9a",x"cf",x"4a"),
   624 => (x"72",x"48",x"c3",x"92"),
   625 => (x"48",x"4a",x"70",x"30"),
   626 => (x"79",x"70",x"b0",x"69"),
   627 => (x"48",x"f4",x"e7",x"c0"),
   628 => (x"e7",x"c0",x"78",x"c0"),
   629 => (x"78",x"c0",x"48",x"f0"),
   630 => (x"49",x"f4",x"cf",x"c1"),
   631 => (x"70",x"87",x"e8",x"fa"),
   632 => (x"aa",x"b7",x"c0",x"4a"),
   633 => (x"87",x"f4",x"fd",x"03"),
   634 => (x"4b",x"26",x"48",x"c0"),
   635 => (x"00",x"00",x"4f",x"26"),
   636 => (x"00",x"00",x"00",x"00"),
   637 => (x"00",x"00",x"00",x"00"),
   638 => (x"72",x"4a",x"c0",x"1e"),
   639 => (x"c0",x"91",x"c4",x"49"),
   640 => (x"c0",x"81",x"cc",x"e9"),
   641 => (x"d0",x"82",x"c1",x"79"),
   642 => (x"ee",x"04",x"aa",x"b7"),
   643 => (x"0e",x"4f",x"26",x"87"),
   644 => (x"5d",x"5c",x"5b",x"5e"),
   645 => (x"f9",x"4d",x"71",x"0e"),
   646 => (x"4a",x"75",x"87",x"dd"),
   647 => (x"92",x"2a",x"b7",x"c4"),
   648 => (x"82",x"cc",x"e9",x"c0"),
   649 => (x"9c",x"cf",x"4c",x"75"),
   650 => (x"49",x"6a",x"94",x"c2"),
   651 => (x"c3",x"2b",x"74",x"4b"),
   652 => (x"74",x"48",x"c2",x"9b"),
   653 => (x"ff",x"4c",x"70",x"30"),
   654 => (x"71",x"48",x"74",x"bc"),
   655 => (x"f8",x"7a",x"70",x"98"),
   656 => (x"48",x"73",x"87",x"ed"),
   657 => (x"4c",x"26",x"4d",x"26"),
   658 => (x"4f",x"26",x"4b",x"26"),
   659 => (x"00",x"00",x"00",x"00"),
   660 => (x"00",x"00",x"00",x"00"),
   661 => (x"00",x"00",x"00",x"00"),
   662 => (x"00",x"00",x"00",x"00"),
   663 => (x"00",x"00",x"00",x"00"),
   664 => (x"00",x"00",x"00",x"00"),
   665 => (x"00",x"00",x"00",x"00"),
   666 => (x"00",x"00",x"00",x"00"),
   667 => (x"00",x"00",x"00",x"00"),
   668 => (x"00",x"00",x"00",x"00"),
   669 => (x"00",x"00",x"00",x"00"),
   670 => (x"00",x"00",x"00",x"00"),
   671 => (x"00",x"00",x"00",x"00"),
   672 => (x"00",x"00",x"00",x"00"),
   673 => (x"00",x"00",x"00",x"00"),
   674 => (x"00",x"00",x"00",x"00"),
   675 => (x"48",x"d0",x"ff",x"1e"),
   676 => (x"71",x"78",x"e1",x"c8"),
   677 => (x"08",x"d4",x"ff",x"48"),
   678 => (x"48",x"66",x"c4",x"78"),
   679 => (x"78",x"08",x"d4",x"ff"),
   680 => (x"71",x"1e",x"4f",x"26"),
   681 => (x"49",x"66",x"c4",x"4a"),
   682 => (x"ff",x"49",x"72",x"1e"),
   683 => (x"d0",x"ff",x"87",x"de"),
   684 => (x"78",x"e0",x"c0",x"48"),
   685 => (x"4f",x"26",x"8e",x"fc"),
   686 => (x"71",x"1e",x"73",x"1e"),
   687 => (x"49",x"66",x"c8",x"4b"),
   688 => (x"c1",x"4a",x"73",x"1e"),
   689 => (x"ff",x"49",x"a2",x"e0"),
   690 => (x"8e",x"fc",x"87",x"d8"),
   691 => (x"4f",x"26",x"4b",x"26"),
   692 => (x"48",x"d0",x"ff",x"1e"),
   693 => (x"71",x"78",x"c9",x"c8"),
   694 => (x"08",x"d4",x"ff",x"48"),
   695 => (x"1e",x"4f",x"26",x"78"),
   696 => (x"eb",x"49",x"4a",x"71"),
   697 => (x"48",x"d0",x"ff",x"87"),
   698 => (x"4f",x"26",x"78",x"c8"),
   699 => (x"71",x"1e",x"73",x"1e"),
   700 => (x"cc",x"d0",x"c1",x"4b"),
   701 => (x"87",x"c3",x"02",x"bf"),
   702 => (x"ff",x"87",x"eb",x"c2"),
   703 => (x"c9",x"c8",x"48",x"d0"),
   704 => (x"c0",x"48",x"73",x"78"),
   705 => (x"d4",x"ff",x"b0",x"e0"),
   706 => (x"d0",x"c1",x"78",x"08"),
   707 => (x"78",x"c0",x"48",x"c0"),
   708 => (x"c5",x"02",x"66",x"c8"),
   709 => (x"49",x"ff",x"c3",x"87"),
   710 => (x"49",x"c0",x"87",x"c2"),
   711 => (x"59",x"c8",x"d0",x"c1"),
   712 => (x"c6",x"02",x"66",x"cc"),
   713 => (x"d5",x"d5",x"c5",x"87"),
   714 => (x"cf",x"87",x"c4",x"4a"),
   715 => (x"c1",x"4a",x"ff",x"ff"),
   716 => (x"c1",x"5a",x"cc",x"d0"),
   717 => (x"c1",x"48",x"cc",x"d0"),
   718 => (x"26",x"4b",x"26",x"78"),
   719 => (x"5b",x"5e",x"0e",x"4f"),
   720 => (x"71",x"0e",x"5d",x"5c"),
   721 => (x"c8",x"d0",x"c1",x"4d"),
   722 => (x"9d",x"75",x"4b",x"bf"),
   723 => (x"49",x"87",x"cb",x"02"),
   724 => (x"eb",x"c0",x"91",x"c8"),
   725 => (x"82",x"71",x"4a",x"e4"),
   726 => (x"ef",x"c0",x"87",x"c4"),
   727 => (x"4c",x"c0",x"4a",x"e4"),
   728 => (x"99",x"73",x"49",x"12"),
   729 => (x"bf",x"c4",x"d0",x"c1"),
   730 => (x"ff",x"b8",x"71",x"48"),
   731 => (x"c1",x"78",x"08",x"d4"),
   732 => (x"c8",x"84",x"2b",x"b7"),
   733 => (x"e7",x"04",x"ac",x"b7"),
   734 => (x"c0",x"d0",x"c1",x"87"),
   735 => (x"80",x"c8",x"48",x"bf"),
   736 => (x"58",x"c4",x"d0",x"c1"),
   737 => (x"4c",x"26",x"4d",x"26"),
   738 => (x"4f",x"26",x"4b",x"26"),
   739 => (x"71",x"1e",x"73",x"1e"),
   740 => (x"9a",x"4a",x"13",x"4b"),
   741 => (x"72",x"87",x"cb",x"02"),
   742 => (x"87",x"e1",x"fe",x"49"),
   743 => (x"05",x"9a",x"4a",x"13"),
   744 => (x"4b",x"26",x"87",x"f5"),
   745 => (x"c1",x"1e",x"4f",x"26"),
   746 => (x"49",x"bf",x"c0",x"d0"),
   747 => (x"48",x"c0",x"d0",x"c1"),
   748 => (x"c4",x"78",x"a1",x"c1"),
   749 => (x"03",x"a9",x"b7",x"c0"),
   750 => (x"d4",x"ff",x"87",x"db"),
   751 => (x"c4",x"d0",x"c1",x"48"),
   752 => (x"d0",x"c1",x"78",x"bf"),
   753 => (x"c1",x"49",x"bf",x"c0"),
   754 => (x"c1",x"48",x"c0",x"d0"),
   755 => (x"c0",x"c4",x"78",x"a1"),
   756 => (x"e5",x"04",x"a9",x"b7"),
   757 => (x"48",x"d0",x"ff",x"87"),
   758 => (x"d0",x"c1",x"78",x"c8"),
   759 => (x"78",x"c0",x"48",x"cc"),
   760 => (x"00",x"00",x"4f",x"26"),
   761 => (x"00",x"00",x"00",x"00"),
   762 => (x"00",x"00",x"00",x"00"),
   763 => (x"5f",x"00",x"00",x"00"),
   764 => (x"00",x"00",x"00",x"5f"),
   765 => (x"00",x"03",x"03",x"00"),
   766 => (x"00",x"00",x"03",x"03"),
   767 => (x"14",x"7f",x"7f",x"14"),
   768 => (x"00",x"14",x"7f",x"7f"),
   769 => (x"6b",x"2e",x"24",x"00"),
   770 => (x"00",x"12",x"3a",x"6b"),
   771 => (x"18",x"36",x"6a",x"4c"),
   772 => (x"00",x"32",x"56",x"6c"),
   773 => (x"59",x"4f",x"7e",x"30"),
   774 => (x"40",x"68",x"3a",x"77"),
   775 => (x"07",x"04",x"00",x"00"),
   776 => (x"00",x"00",x"00",x"03"),
   777 => (x"3e",x"1c",x"00",x"00"),
   778 => (x"00",x"00",x"41",x"63"),
   779 => (x"63",x"41",x"00",x"00"),
   780 => (x"00",x"00",x"1c",x"3e"),
   781 => (x"1c",x"3e",x"2a",x"08"),
   782 => (x"08",x"2a",x"3e",x"1c"),
   783 => (x"3e",x"08",x"08",x"00"),
   784 => (x"00",x"08",x"08",x"3e"),
   785 => (x"e0",x"80",x"00",x"00"),
   786 => (x"00",x"00",x"00",x"60"),
   787 => (x"08",x"08",x"08",x"00"),
   788 => (x"00",x"08",x"08",x"08"),
   789 => (x"60",x"00",x"00",x"00"),
   790 => (x"00",x"00",x"00",x"60"),
   791 => (x"18",x"30",x"60",x"40"),
   792 => (x"01",x"03",x"06",x"0c"),
   793 => (x"59",x"7f",x"3e",x"00"),
   794 => (x"00",x"3e",x"7f",x"4d"),
   795 => (x"7f",x"06",x"04",x"00"),
   796 => (x"00",x"00",x"00",x"7f"),
   797 => (x"71",x"63",x"42",x"00"),
   798 => (x"00",x"46",x"4f",x"59"),
   799 => (x"49",x"63",x"22",x"00"),
   800 => (x"00",x"36",x"7f",x"49"),
   801 => (x"13",x"16",x"1c",x"18"),
   802 => (x"00",x"10",x"7f",x"7f"),
   803 => (x"45",x"67",x"27",x"00"),
   804 => (x"00",x"39",x"7d",x"45"),
   805 => (x"4b",x"7e",x"3c",x"00"),
   806 => (x"00",x"30",x"79",x"49"),
   807 => (x"71",x"01",x"01",x"00"),
   808 => (x"00",x"07",x"0f",x"79"),
   809 => (x"49",x"7f",x"36",x"00"),
   810 => (x"00",x"36",x"7f",x"49"),
   811 => (x"49",x"4f",x"06",x"00"),
   812 => (x"00",x"1e",x"3f",x"69"),
   813 => (x"66",x"00",x"00",x"00"),
   814 => (x"00",x"00",x"00",x"66"),
   815 => (x"e6",x"80",x"00",x"00"),
   816 => (x"00",x"00",x"00",x"66"),
   817 => (x"14",x"08",x"08",x"00"),
   818 => (x"00",x"22",x"22",x"14"),
   819 => (x"14",x"14",x"14",x"00"),
   820 => (x"00",x"14",x"14",x"14"),
   821 => (x"14",x"22",x"22",x"00"),
   822 => (x"00",x"08",x"08",x"14"),
   823 => (x"51",x"03",x"02",x"00"),
   824 => (x"00",x"06",x"0f",x"59"),
   825 => (x"5d",x"41",x"7f",x"3e"),
   826 => (x"00",x"1e",x"1f",x"55"),
   827 => (x"09",x"7f",x"7e",x"00"),
   828 => (x"00",x"7e",x"7f",x"09"),
   829 => (x"49",x"7f",x"7f",x"00"),
   830 => (x"00",x"36",x"7f",x"49"),
   831 => (x"63",x"3e",x"1c",x"00"),
   832 => (x"00",x"41",x"41",x"41"),
   833 => (x"41",x"7f",x"7f",x"00"),
   834 => (x"00",x"1c",x"3e",x"63"),
   835 => (x"49",x"7f",x"7f",x"00"),
   836 => (x"00",x"41",x"41",x"49"),
   837 => (x"09",x"7f",x"7f",x"00"),
   838 => (x"00",x"01",x"01",x"09"),
   839 => (x"41",x"7f",x"3e",x"00"),
   840 => (x"00",x"7a",x"7b",x"49"),
   841 => (x"08",x"7f",x"7f",x"00"),
   842 => (x"00",x"7f",x"7f",x"08"),
   843 => (x"7f",x"41",x"00",x"00"),
   844 => (x"00",x"00",x"41",x"7f"),
   845 => (x"40",x"60",x"20",x"00"),
   846 => (x"00",x"3f",x"7f",x"40"),
   847 => (x"1c",x"08",x"7f",x"7f"),
   848 => (x"00",x"41",x"63",x"36"),
   849 => (x"40",x"7f",x"7f",x"00"),
   850 => (x"00",x"40",x"40",x"40"),
   851 => (x"0c",x"06",x"7f",x"7f"),
   852 => (x"00",x"7f",x"7f",x"06"),
   853 => (x"0c",x"06",x"7f",x"7f"),
   854 => (x"00",x"7f",x"7f",x"18"),
   855 => (x"41",x"7f",x"3e",x"00"),
   856 => (x"00",x"3e",x"7f",x"41"),
   857 => (x"09",x"7f",x"7f",x"00"),
   858 => (x"00",x"06",x"0f",x"09"),
   859 => (x"61",x"41",x"7f",x"3e"),
   860 => (x"00",x"40",x"7e",x"7f"),
   861 => (x"09",x"7f",x"7f",x"00"),
   862 => (x"00",x"66",x"7f",x"19"),
   863 => (x"4d",x"6f",x"26",x"00"),
   864 => (x"00",x"32",x"7b",x"59"),
   865 => (x"7f",x"01",x"01",x"00"),
   866 => (x"00",x"01",x"01",x"7f"),
   867 => (x"40",x"7f",x"3f",x"00"),
   868 => (x"00",x"3f",x"7f",x"40"),
   869 => (x"70",x"3f",x"0f",x"00"),
   870 => (x"00",x"0f",x"3f",x"70"),
   871 => (x"18",x"30",x"7f",x"7f"),
   872 => (x"00",x"7f",x"7f",x"30"),
   873 => (x"1c",x"36",x"63",x"41"),
   874 => (x"41",x"63",x"36",x"1c"),
   875 => (x"7c",x"06",x"03",x"01"),
   876 => (x"01",x"03",x"06",x"7c"),
   877 => (x"4d",x"59",x"71",x"61"),
   878 => (x"00",x"41",x"43",x"47"),
   879 => (x"7f",x"7f",x"00",x"00"),
   880 => (x"00",x"00",x"41",x"41"),
   881 => (x"0c",x"06",x"03",x"01"),
   882 => (x"40",x"60",x"30",x"18"),
   883 => (x"41",x"41",x"00",x"00"),
   884 => (x"00",x"00",x"7f",x"7f"),
   885 => (x"03",x"06",x"0c",x"08"),
   886 => (x"00",x"08",x"0c",x"06"),
   887 => (x"80",x"80",x"80",x"80"),
   888 => (x"00",x"80",x"80",x"80"),
   889 => (x"03",x"00",x"00",x"00"),
   890 => (x"00",x"00",x"04",x"07"),
   891 => (x"54",x"74",x"20",x"00"),
   892 => (x"00",x"78",x"7c",x"54"),
   893 => (x"44",x"7f",x"7f",x"00"),
   894 => (x"00",x"38",x"7c",x"44"),
   895 => (x"44",x"7c",x"38",x"00"),
   896 => (x"00",x"00",x"44",x"44"),
   897 => (x"44",x"7c",x"38",x"00"),
   898 => (x"00",x"7f",x"7f",x"44"),
   899 => (x"54",x"7c",x"38",x"00"),
   900 => (x"00",x"18",x"5c",x"54"),
   901 => (x"7f",x"7e",x"04",x"00"),
   902 => (x"00",x"00",x"05",x"05"),
   903 => (x"a4",x"bc",x"18",x"00"),
   904 => (x"00",x"7c",x"fc",x"a4"),
   905 => (x"04",x"7f",x"7f",x"00"),
   906 => (x"00",x"78",x"7c",x"04"),
   907 => (x"3d",x"00",x"00",x"00"),
   908 => (x"00",x"00",x"40",x"7d"),
   909 => (x"80",x"80",x"80",x"00"),
   910 => (x"00",x"00",x"7d",x"fd"),
   911 => (x"10",x"7f",x"7f",x"00"),
   912 => (x"00",x"44",x"6c",x"38"),
   913 => (x"3f",x"00",x"00",x"00"),
   914 => (x"00",x"00",x"40",x"7f"),
   915 => (x"18",x"0c",x"7c",x"7c"),
   916 => (x"00",x"78",x"7c",x"0c"),
   917 => (x"04",x"7c",x"7c",x"00"),
   918 => (x"00",x"78",x"7c",x"04"),
   919 => (x"44",x"7c",x"38",x"00"),
   920 => (x"00",x"38",x"7c",x"44"),
   921 => (x"24",x"fc",x"fc",x"00"),
   922 => (x"00",x"18",x"3c",x"24"),
   923 => (x"24",x"3c",x"18",x"00"),
   924 => (x"00",x"fc",x"fc",x"24"),
   925 => (x"04",x"7c",x"7c",x"00"),
   926 => (x"00",x"08",x"0c",x"04"),
   927 => (x"54",x"5c",x"48",x"00"),
   928 => (x"00",x"20",x"74",x"54"),
   929 => (x"7f",x"3f",x"04",x"00"),
   930 => (x"00",x"00",x"44",x"44"),
   931 => (x"40",x"7c",x"3c",x"00"),
   932 => (x"00",x"7c",x"7c",x"40"),
   933 => (x"60",x"3c",x"1c",x"00"),
   934 => (x"00",x"1c",x"3c",x"60"),
   935 => (x"30",x"60",x"7c",x"3c"),
   936 => (x"00",x"3c",x"7c",x"60"),
   937 => (x"10",x"38",x"6c",x"44"),
   938 => (x"00",x"44",x"6c",x"38"),
   939 => (x"e0",x"bc",x"1c",x"00"),
   940 => (x"00",x"1c",x"3c",x"60"),
   941 => (x"74",x"64",x"44",x"00"),
   942 => (x"00",x"44",x"4c",x"5c"),
   943 => (x"3e",x"08",x"08",x"00"),
   944 => (x"00",x"41",x"41",x"77"),
   945 => (x"7f",x"00",x"00",x"00"),
   946 => (x"00",x"00",x"00",x"7f"),
   947 => (x"77",x"41",x"41",x"00"),
   948 => (x"00",x"08",x"08",x"3e"),
   949 => (x"03",x"01",x"01",x"02"),
   950 => (x"00",x"01",x"02",x"02"),
   951 => (x"7f",x"7f",x"7f",x"7f"),
   952 => (x"00",x"7f",x"7f",x"7f"),
   953 => (x"1c",x"1c",x"08",x"08"),
   954 => (x"7f",x"7f",x"3e",x"3e"),
   955 => (x"3e",x"3e",x"7f",x"7f"),
   956 => (x"08",x"08",x"1c",x"1c"),
   957 => (x"7c",x"18",x"10",x"00"),
   958 => (x"00",x"10",x"18",x"7c"),
   959 => (x"7c",x"30",x"10",x"00"),
   960 => (x"00",x"10",x"30",x"7c"),
   961 => (x"60",x"60",x"30",x"10"),
   962 => (x"00",x"06",x"1e",x"78"),
   963 => (x"18",x"3c",x"66",x"42"),
   964 => (x"00",x"42",x"66",x"3c"),
   965 => (x"c2",x"6a",x"38",x"78"),
   966 => (x"00",x"38",x"6c",x"c6"),
   967 => (x"60",x"00",x"00",x"60"),
   968 => (x"00",x"60",x"00",x"00"),
   969 => (x"5c",x"5b",x"5e",x"0e"),
   970 => (x"86",x"fc",x"0e",x"5d"),
   971 => (x"d0",x"c1",x"7e",x"71"),
   972 => (x"c0",x"4c",x"bf",x"d4"),
   973 => (x"c4",x"1e",x"c0",x"4b"),
   974 => (x"c4",x"02",x"ab",x"66"),
   975 => (x"c2",x"4d",x"c0",x"87"),
   976 => (x"75",x"4d",x"c1",x"87"),
   977 => (x"ee",x"49",x"73",x"1e"),
   978 => (x"86",x"c8",x"87",x"e2"),
   979 => (x"ef",x"49",x"e0",x"c0"),
   980 => (x"a4",x"c4",x"87",x"eb"),
   981 => (x"f0",x"49",x"6a",x"4a"),
   982 => (x"c9",x"f1",x"87",x"f2"),
   983 => (x"c1",x"84",x"cc",x"87"),
   984 => (x"ab",x"b7",x"c8",x"83"),
   985 => (x"87",x"cd",x"ff",x"04"),
   986 => (x"4d",x"26",x"8e",x"fc"),
   987 => (x"4b",x"26",x"4c",x"26"),
   988 => (x"71",x"1e",x"4f",x"26"),
   989 => (x"d8",x"d0",x"c1",x"4a"),
   990 => (x"d8",x"d0",x"c1",x"5a"),
   991 => (x"49",x"78",x"c7",x"48"),
   992 => (x"26",x"87",x"e1",x"fe"),
   993 => (x"1e",x"73",x"1e",x"4f"),
   994 => (x"b7",x"c0",x"4a",x"71"),
   995 => (x"87",x"d3",x"03",x"aa"),
   996 => (x"bf",x"e0",x"cb",x"c1"),
   997 => (x"c1",x"87",x"c4",x"05"),
   998 => (x"c0",x"87",x"c2",x"4b"),
   999 => (x"e4",x"cb",x"c1",x"4b"),
  1000 => (x"c1",x"87",x"c4",x"5b"),
  1001 => (x"fc",x"5a",x"e4",x"cb"),
  1002 => (x"e0",x"cb",x"c1",x"48"),
  1003 => (x"c1",x"4a",x"78",x"bf"),
  1004 => (x"a2",x"c0",x"c1",x"9a"),
  1005 => (x"87",x"e7",x"ec",x"49"),
  1006 => (x"4f",x"26",x"4b",x"26"),
  1007 => (x"c4",x"4a",x"71",x"1e"),
  1008 => (x"49",x"72",x"1e",x"66"),
  1009 => (x"fc",x"87",x"f1",x"eb"),
  1010 => (x"1e",x"4f",x"26",x"8e"),
  1011 => (x"c3",x"48",x"d4",x"ff"),
  1012 => (x"d0",x"ff",x"78",x"ff"),
  1013 => (x"78",x"e1",x"c0",x"48"),
  1014 => (x"c1",x"48",x"d4",x"ff"),
  1015 => (x"c4",x"48",x"71",x"78"),
  1016 => (x"08",x"d4",x"ff",x"30"),
  1017 => (x"48",x"d0",x"ff",x"78"),
  1018 => (x"26",x"78",x"e0",x"c0"),
  1019 => (x"5b",x"5e",x"0e",x"4f"),
  1020 => (x"ec",x"0e",x"5d",x"5c"),
  1021 => (x"48",x"a6",x"c8",x"86"),
  1022 => (x"c4",x"7e",x"78",x"c0"),
  1023 => (x"78",x"bf",x"ec",x"80"),
  1024 => (x"d0",x"c1",x"80",x"f8"),
  1025 => (x"e8",x"78",x"bf",x"d4"),
  1026 => (x"cb",x"c1",x"4c",x"bf"),
  1027 => (x"e4",x"49",x"bf",x"e0"),
  1028 => (x"ee",x"cb",x"87",x"f7"),
  1029 => (x"87",x"cc",x"cb",x"49"),
  1030 => (x"c7",x"58",x"a6",x"d4"),
  1031 => (x"87",x"ef",x"e7",x"49"),
  1032 => (x"c9",x"05",x"98",x"70"),
  1033 => (x"49",x"66",x"cc",x"87"),
  1034 => (x"c1",x"02",x"99",x"c1"),
  1035 => (x"66",x"d0",x"87",x"c4"),
  1036 => (x"ec",x"7e",x"c1",x"4d"),
  1037 => (x"cb",x"c1",x"4b",x"bf"),
  1038 => (x"e4",x"49",x"bf",x"e0"),
  1039 => (x"49",x"75",x"87",x"cb"),
  1040 => (x"70",x"87",x"ed",x"ca"),
  1041 => (x"87",x"d7",x"02",x"98"),
  1042 => (x"bf",x"c8",x"cb",x"c1"),
  1043 => (x"c1",x"b9",x"c1",x"49"),
  1044 => (x"71",x"59",x"cc",x"cb"),
  1045 => (x"cb",x"87",x"f4",x"fd"),
  1046 => (x"c7",x"ca",x"49",x"ee"),
  1047 => (x"c7",x"4d",x"70",x"87"),
  1048 => (x"87",x"eb",x"e6",x"49"),
  1049 => (x"ff",x"05",x"98",x"70"),
  1050 => (x"49",x"73",x"87",x"c7"),
  1051 => (x"fe",x"05",x"99",x"c1"),
  1052 => (x"02",x"6e",x"87",x"ff"),
  1053 => (x"c1",x"87",x"e3",x"c0"),
  1054 => (x"4a",x"bf",x"e0",x"cb"),
  1055 => (x"cb",x"c1",x"ba",x"c1"),
  1056 => (x"0a",x"fc",x"5a",x"e4"),
  1057 => (x"9a",x"c1",x"0a",x"7a"),
  1058 => (x"49",x"a2",x"c0",x"c1"),
  1059 => (x"c1",x"87",x"d0",x"e9"),
  1060 => (x"fa",x"e5",x"49",x"da"),
  1061 => (x"48",x"a6",x"c8",x"87"),
  1062 => (x"cb",x"c1",x"78",x"c1"),
  1063 => (x"c1",x"05",x"bf",x"e0"),
  1064 => (x"c0",x"c8",x"87",x"c5"),
  1065 => (x"cb",x"c1",x"4d",x"c0"),
  1066 => (x"49",x"13",x"4b",x"cc"),
  1067 => (x"87",x"df",x"e5",x"49"),
  1068 => (x"c2",x"02",x"98",x"70"),
  1069 => (x"c1",x"b4",x"75",x"87"),
  1070 => (x"ff",x"05",x"2d",x"b7"),
  1071 => (x"49",x"74",x"87",x"ec"),
  1072 => (x"71",x"99",x"ff",x"c3"),
  1073 => (x"fb",x"49",x"c0",x"1e"),
  1074 => (x"49",x"74",x"87",x"f2"),
  1075 => (x"71",x"29",x"b7",x"c8"),
  1076 => (x"fb",x"49",x"c1",x"1e"),
  1077 => (x"86",x"c8",x"87",x"e6"),
  1078 => (x"e4",x"49",x"fd",x"c3"),
  1079 => (x"fa",x"c3",x"87",x"f1"),
  1080 => (x"87",x"eb",x"e4",x"49"),
  1081 => (x"74",x"87",x"d4",x"c7"),
  1082 => (x"99",x"ff",x"c3",x"49"),
  1083 => (x"71",x"2c",x"b7",x"c8"),
  1084 => (x"02",x"9c",x"74",x"b4"),
  1085 => (x"cb",x"c1",x"87",x"df"),
  1086 => (x"c7",x"49",x"bf",x"dc"),
  1087 => (x"98",x"70",x"87",x"f2"),
  1088 => (x"87",x"c4",x"c0",x"05"),
  1089 => (x"87",x"d3",x"4c",x"c0"),
  1090 => (x"c7",x"49",x"e0",x"c2"),
  1091 => (x"cb",x"c1",x"87",x"d6"),
  1092 => (x"c6",x"c0",x"58",x"e0"),
  1093 => (x"dc",x"cb",x"c1",x"87"),
  1094 => (x"74",x"78",x"c0",x"48"),
  1095 => (x"05",x"99",x"c8",x"49"),
  1096 => (x"c3",x"87",x"ce",x"c0"),
  1097 => (x"e6",x"e3",x"49",x"f5"),
  1098 => (x"c2",x"49",x"70",x"87"),
  1099 => (x"e7",x"c0",x"02",x"99"),
  1100 => (x"d8",x"d0",x"c1",x"87"),
  1101 => (x"ca",x"c0",x"02",x"bf"),
  1102 => (x"88",x"c1",x"48",x"87"),
  1103 => (x"58",x"dc",x"d0",x"c1"),
  1104 => (x"c4",x"87",x"d0",x"c0"),
  1105 => (x"e0",x"c1",x"4a",x"66"),
  1106 => (x"c0",x"02",x"6a",x"82"),
  1107 => (x"ff",x"4b",x"87",x"c5"),
  1108 => (x"c8",x"0f",x"73",x"49"),
  1109 => (x"78",x"c1",x"48",x"a6"),
  1110 => (x"99",x"c4",x"49",x"74"),
  1111 => (x"87",x"ce",x"c0",x"05"),
  1112 => (x"e2",x"49",x"f2",x"c3"),
  1113 => (x"49",x"70",x"87",x"e9"),
  1114 => (x"c0",x"02",x"99",x"c2"),
  1115 => (x"d0",x"c1",x"87",x"f0"),
  1116 => (x"48",x"7e",x"bf",x"d8"),
  1117 => (x"03",x"a8",x"b7",x"c7"),
  1118 => (x"6e",x"87",x"cb",x"c0"),
  1119 => (x"c1",x"80",x"c1",x"48"),
  1120 => (x"c0",x"58",x"dc",x"d0"),
  1121 => (x"66",x"c4",x"87",x"d3"),
  1122 => (x"80",x"e0",x"c1",x"48"),
  1123 => (x"bf",x"6e",x"7e",x"70"),
  1124 => (x"87",x"c5",x"c0",x"02"),
  1125 => (x"73",x"49",x"fe",x"4b"),
  1126 => (x"48",x"a6",x"c8",x"0f"),
  1127 => (x"fd",x"c3",x"78",x"c1"),
  1128 => (x"87",x"eb",x"e1",x"49"),
  1129 => (x"99",x"c2",x"49",x"70"),
  1130 => (x"87",x"e9",x"c0",x"02"),
  1131 => (x"bf",x"d8",x"d0",x"c1"),
  1132 => (x"87",x"c9",x"c0",x"02"),
  1133 => (x"48",x"d8",x"d0",x"c1"),
  1134 => (x"d3",x"c0",x"78",x"c0"),
  1135 => (x"48",x"66",x"c4",x"87"),
  1136 => (x"70",x"80",x"e0",x"c1"),
  1137 => (x"02",x"bf",x"6e",x"7e"),
  1138 => (x"4b",x"87",x"c5",x"c0"),
  1139 => (x"0f",x"73",x"49",x"fd"),
  1140 => (x"c1",x"48",x"a6",x"c8"),
  1141 => (x"49",x"fa",x"c3",x"78"),
  1142 => (x"70",x"87",x"f4",x"e0"),
  1143 => (x"02",x"99",x"c2",x"49"),
  1144 => (x"c1",x"87",x"ed",x"c0"),
  1145 => (x"48",x"bf",x"d8",x"d0"),
  1146 => (x"03",x"a8",x"b7",x"c7"),
  1147 => (x"c1",x"87",x"c9",x"c0"),
  1148 => (x"c7",x"48",x"d8",x"d0"),
  1149 => (x"87",x"d3",x"c0",x"78"),
  1150 => (x"c1",x"48",x"66",x"c4"),
  1151 => (x"7e",x"70",x"80",x"e0"),
  1152 => (x"c0",x"02",x"bf",x"6e"),
  1153 => (x"fc",x"4b",x"87",x"c5"),
  1154 => (x"c8",x"0f",x"73",x"49"),
  1155 => (x"78",x"c1",x"48",x"a6"),
  1156 => (x"d0",x"c1",x"7e",x"c0"),
  1157 => (x"50",x"c0",x"48",x"d0"),
  1158 => (x"c3",x"49",x"ee",x"cb"),
  1159 => (x"a6",x"d4",x"87",x"c6"),
  1160 => (x"d0",x"d0",x"c1",x"58"),
  1161 => (x"c1",x"05",x"bf",x"97"),
  1162 => (x"49",x"74",x"87",x"de"),
  1163 => (x"05",x"99",x"f0",x"c3"),
  1164 => (x"c1",x"87",x"cd",x"c0"),
  1165 => (x"df",x"ff",x"49",x"da"),
  1166 => (x"98",x"70",x"87",x"d5"),
  1167 => (x"87",x"c8",x"c1",x"02"),
  1168 => (x"bf",x"e8",x"7e",x"c1"),
  1169 => (x"ff",x"c3",x"49",x"4b"),
  1170 => (x"2b",x"b7",x"c8",x"99"),
  1171 => (x"cb",x"c1",x"b3",x"71"),
  1172 => (x"ff",x"49",x"bf",x"e0"),
  1173 => (x"d0",x"87",x"f2",x"db"),
  1174 => (x"d3",x"c2",x"49",x"66"),
  1175 => (x"02",x"98",x"70",x"87"),
  1176 => (x"c1",x"87",x"c6",x"c0"),
  1177 => (x"c1",x"48",x"d0",x"d0"),
  1178 => (x"d0",x"d0",x"c1",x"50"),
  1179 => (x"c0",x"05",x"bf",x"97"),
  1180 => (x"49",x"73",x"87",x"d6"),
  1181 => (x"05",x"99",x"f0",x"c3"),
  1182 => (x"c1",x"87",x"c5",x"ff"),
  1183 => (x"de",x"ff",x"49",x"da"),
  1184 => (x"98",x"70",x"87",x"cd"),
  1185 => (x"87",x"f8",x"fe",x"05"),
  1186 => (x"e0",x"c0",x"02",x"6e"),
  1187 => (x"48",x"a6",x"cc",x"87"),
  1188 => (x"bf",x"d8",x"d0",x"c1"),
  1189 => (x"49",x"66",x"cc",x"78"),
  1190 => (x"66",x"c4",x"91",x"cc"),
  1191 => (x"70",x"80",x"71",x"48"),
  1192 => (x"02",x"bf",x"6e",x"7e"),
  1193 => (x"4b",x"87",x"c6",x"c0"),
  1194 => (x"73",x"49",x"66",x"cc"),
  1195 => (x"02",x"66",x"c8",x"0f"),
  1196 => (x"c1",x"87",x"c8",x"c0"),
  1197 => (x"49",x"bf",x"d8",x"d0"),
  1198 => (x"ec",x"87",x"e9",x"f1"),
  1199 => (x"26",x"4d",x"26",x"8e"),
  1200 => (x"26",x"4b",x"26",x"4c"),
  1201 => (x"00",x"00",x"00",x"4f"),
  1202 => (x"00",x"00",x"00",x"00"),
  1203 => (x"14",x"11",x"12",x"58"),
  1204 => (x"23",x"1c",x"1b",x"1d"),
  1205 => (x"94",x"91",x"59",x"5a"),
  1206 => (x"f4",x"eb",x"f2",x"f5"),
  1207 => (x"00",x"00",x"00",x"00"),
  1208 => (x"00",x"00",x"00",x"00"),
  1209 => (x"ff",x"4a",x"71",x"1e"),
  1210 => (x"72",x"49",x"bf",x"c8"),
  1211 => (x"4f",x"26",x"48",x"a1"),
  1212 => (x"bf",x"c8",x"ff",x"1e"),
  1213 => (x"c0",x"c0",x"fe",x"89"),
  1214 => (x"a9",x"c0",x"c0",x"c0"),
  1215 => (x"c0",x"87",x"c4",x"01"),
  1216 => (x"c1",x"87",x"c2",x"4a"),
  1217 => (x"26",x"48",x"72",x"4a"),
  1218 => (x"00",x"08",x"5f",x"4f"),
  1219 => (x"00",x"08",x"5f",x"00"),
		others => (others => x"00")
	);
	signal q1_local : word_t;

	-- Altera Quartus attributes
	attribute ramstyle: string;
	attribute ramstyle of ram: signal is "no_rw_check";

begin  -- rtl

	addr1 <= to_integer(unsigned(addr(ADDR_WIDTH-1 downto 0)));

	-- Reorganize the read data from the RAM to match the output
	q(7 downto 0) <= q1_local(3);
	q(15 downto 8) <= q1_local(2);
	q(23 downto 16) <= q1_local(1);
	q(31 downto 24) <= q1_local(0);

	process(clk)
	begin
		if(rising_edge(clk)) then 
			if(we = '1') then
				-- edit this code if using other than four bytes per word
				if (bytesel(3) = '1') then
					ram(addr1)(3) <= d(7 downto 0);
				end if;
				if (bytesel(2) = '1') then
					ram(addr1)(2) <= d(15 downto 8);
				end if;
				if (bytesel(1) = '1') then
					ram(addr1)(1) <= d(23 downto 16);
				end if;
				if (bytesel(0) = '1') then
					ram(addr1)(0) <= d(31 downto 24);
				end if;
			end if;
			q1_local <= ram(addr1);
		end if;
	end process;
  
end rtl;

